module shift_reg(reg_out, reg_in, clock);

output [3:0] reg_out;
input [3:0] reg_in;
input clock;

//internals not shown

endmodule
