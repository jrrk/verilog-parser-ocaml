
module hello_top;

initial
	$hello_verilog; //Invoke the user defined task $hello_verilog

endmodule


